module pre_input_transposer #(
    parameter DATA_WIDTH    = 39
)
(
    input   wire    clk,
    input   wire    rst_n,

    input   wire                        i_ibuf_reset,
    output  wire                        o_ibuf_done,

    input   wire                        i_ibuf_wren,
    input   wire    [11:0]              i_ibuf_addr,    // 0 ~ 3071
    input   wire    [2*DATA_WIDTH-1:0]  i_ibuf_data,

    output  wire    [47:0]              o_ibuf_wren,    // p5b7 ~ p0b7 ~ p0b0 : p = polyn, b = bank = 1/8 polyn
    output  wire    [71:0]              o_ibuf_addr,    // 9 * 8
    output  wire    [8*DATA_WIDTH-1:0]  o_ibuf_data     // 35/39 * 8
);


    reg input_completed_r;
    wire input_completed;       // all 8 polynomials received
    wire output_completed;      // all 8 polynomials saved to ram
    assign o_ibuf_done = input_completed_r & output_completed;
    

    /* input logic begin */
    wire [10:0] count_i_coeff;   // number of coeff in a polynomial received
    wire [2:0] count_i_polyn;   // number of polyn received

    assign count_i_coeff = i_ibuf_addr[10:0];
    assign count_i_polyn = i_ibuf_addr[11:9];
    assign input_completed = (i_ibuf_addr == 12'h7ff);

    always @ (posedge clk or negedge rst_n) begin
        if (~rst_n)
            input_completed_r <= 1'b0;
        else if (i_ibuf_reset)
            input_completed_r <= 1'b0;
        else if (o_ibuf_done)
            input_completed_r <= 1'b0;
        else if (input_completed)
            input_completed_r <= 1'b1;
        else
            input_completed_r <= input_completed_r;
    end
    /* input logic end */


    reg [7:0] o_comp;
    assign output_completed = &o_comp[7:0];

    genvar i, j;
    generate
        for (i = 0; i < 8; i = i + 1) begin : gen_buf

            wire iwren;
            wire [7:0] iaddr;
            assign iwren = (count_i_coeff[10:8] == i) && i_ibuf_wren;
            assign iaddr = count_i_coeff[7:0];

            reg [5:0] owren;
            reg [5:0] owren_m1; // lutram delay = 1 cycle
            wire [8:0] oaddr;
            reg [8:0] oaddr_m1; // lutram delay = 1 cycle
            reg [DATA_WIDTH-1:0] odata;

            assign o_ibuf_wren[i*6 +: 6] = owren_m1;
            assign o_ibuf_addr[i*9 +: 9] = oaddr_m1;
            assign o_ibuf_data[i*DATA_WIDTH +: DATA_WIDTH] = odata;

            always @ (posedge clk) begin
                oaddr_m1 <= oaddr;
                owren_m1 <= owren;
            end

            /* instantiate buffer begin */
            wire [2*DATA_WIDTH-1:0] ram_dout;
            wire [2*DATA_WIDTH-1:0] ram_din;
            assign ram_din = i_ibuf_data;

            /*
            xpm_memory_sdpram #(
                .ADDR_WIDTH_A           ( 8                     ),
                .ADDR_WIDTH_B           ( 8                     ),
                .AUTO_SLEEP_TIME        ( 0                     ),
                .BYTE_WRITE_WIDTH_A     ( 2 * DATA_WIDTH        ),
                .CASCADE_HEIGHT         ( 0                     ),
                .CLOCKING_MODE          ( "common_clock"        ),
                .ECC_MODE               ( "no_ecc"              ),
                .MEMORY_INIT_FILE       ( "none"                ),
                .MEMORY_INIT_PARAM      ( "0"                   ),
                .MEMORY_OPTIMIZATION    ( "true"                ),
                .MEMORY_PRIMITIVE       ( "distributed"         ),
                .MEMORY_SIZE            ( 2 * DATA_WIDTH * 256   ),
                .MESSAGE_CONTROL        ( 0                     ),
                .READ_DATA_WIDTH_B      ( 2 * DATA_WIDTH        ),
                .READ_LATENCY_B         ( 1                     ),
                .READ_RESET_VALUE_B     ( "0"                   ),
                .RST_MODE_A             ( "SYNC"                ),
                .RST_MODE_B             ( "SYNC"                ),
                .SIM_ASSERT_CHK         ( 0                     ),
                .USE_EMBEDDED_CONSTRAINT( 0                     ),
                .USE_MEM_INIT           ( 0                     ),
                .WAKEUP_TIME            ( "disable_sleep"       ),
                .WRITE_DATA_WIDTH_A     ( 2 * DATA_WIDTH        ),
                .WRITE_MODE_B           ( "read_first"          )
            )
            i_ibuf_lutram_sdpram (
                .clka   ( clk               ),
                .clkb   ( clk               ),
                .ena    ( 1'b1              ),
                .enb    ( 1'b1              ),
                .addra  ( iaddr[7:0]        ),
                .addrb  ( oaddr[8:1]        ),
                .wea    ( iwren             ),
                .dina   ( ram_din           ),
                .doutb  ( ram_dout          ),
                .regceb ( 1'b1              ),
                .rstb   ( 1'b0              )
            );
            */
            
            sdpram #(
                .ADDR_WIDTH_A        (8),
                .ADDR_WIDTH_B        (8),
                .WRITE_DATA_WIDTH_A  (2 * DATA_WIDTH),
                .READ_DATA_WIDTH_B   (2 * DATA_WIDTH),
                .READ_LATENCY_B      (1),
                .WRITE_MODE_B        (0)  // 0 = read_first
            ) i_ibuf_lutram_sdpram (
                .clka    ( clk               ),
                .clkb    ( clk               ),
                .ena     ( 1'b1              ),
                .enb     ( 1'b1              ),
                .addra   ( iaddr[7:0]        ),
                .addrb   ( oaddr[8:1]        ),
                .wea     ( iwren             ),
                .dina    ( ram_din           ),
                .doutb   ( ram_dout          ),
                .regceb  ( 1'b1              ),
                .rstb    ( 1'b0              )
            );

            always @ (*) begin
                odata = 'b0;
                case (oaddr_m1[0])
                    1'd0: odata = ram_dout[0 * DATA_WIDTH +: DATA_WIDTH];
                    1'd1: odata = ram_dout[1 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd2: odata = ram_dout[2 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd3: odata = ram_dout[3 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd4: odata = ram_dout[4 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd5: odata = ram_dout[5 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd6: odata = ram_dout[6 * DATA_WIDTH +: DATA_WIDTH];
                    //3'd7: odata = ram_dout[7 * DATA_WIDTH +: DATA_WIDTH];
                endcase
            end
            /* instantiate buffer end */


            /* output logic begin */
            reg vld;
            wire [10:0] count_o_coeff;
            wire [2:0] count_o_polyn;

            assign oaddr = count_o_coeff;

            always @ (posedge clk or negedge rst_n) begin
                if (~rst_n)
                    vld <= 1'b0;
                else if (i_ibuf_reset)
                    vld <= 1'b0;
                else if (count_i_coeff[10:8] == i &&
                         count_i_coeff[5:0] == 6'd62 && // early start
                         i_ibuf_wren)
                    vld <= 1'b1;
                else if (vld && count_o_coeff[10:0] == 11'd2047) // 2047 because we need to count to the max coefficient
                    vld <= 1'b0;
                else
                    vld <= vld;
            end

            counter #(.C_WIDTH(14), . MAX_COUNT('h7FF), .C_INIT(14'd0))
            i_cntr_output(
                .clk        ( clk                               ),
                .clken      ( 1'b1                              ),
                .rst        ( ~rst_n                            ),
                .load       ( i_ibuf_reset                      ),
                .incr       ( vld                               ),
                .decr       ( 1'b0                              ),
                .load_value ( 14'd0                             ),
                .count      ( {count_o_polyn, count_o_coeff}    ),
                .is_zero    (                                   )
            );

            always @ (*) begin
                owren = 'b0;
                if (vld) begin
                    case ({count_o_polyn[0], count_o_coeff[10:9]})
                        3'd0: owren = 6'b00_0001;
                        3'd1: owren = 6'b00_0010;
                        3'd2: owren = 6'b00_0100;
                        3'd3: owren = 6'b00_1000;
                        3'd4: owren = 6'b01_0000;
                        3'd5: owren = 6'b10_0000;
                    endcase
                end
            end
            
            always @ (posedge clk or negedge rst_n) begin
                if (~rst_n)
                    o_comp[i] <= 1'b0;
                else if (i_ibuf_reset)
                    o_comp[i] <= 1'b0;
                else if (o_ibuf_done)
                    o_comp[i] <= 1'b0;
                else if (count_o_coeff == 11'h7FF)
                    o_comp[i] <= 1'b1;
                else
                    o_comp[i] <= o_comp[i];
            end
            /* output logic end */

        end
    endgenerate

endmodule


// Vendor-agnostic simple dual-port RAM (common or independent clocks)
// Port A: write; Port B: read; READ_MODE_B: "read_first"; READ_LATENCY_B >= 1
module sdpram #(
  parameter integer ADDR_WIDTH_A        = 8,
  parameter integer ADDR_WIDTH_B        = 8,
  parameter integer WRITE_DATA_WIDTH_A  = 64,
  parameter integer READ_DATA_WIDTH_B   = 64,
  parameter integer READ_LATENCY_B      = 1,  // >=1
  parameter integer WRITE_MODE_B        = 0   // 0=read_first (modeled)
)(
  input  wire                          clka,
  input  wire                          clkb,
  input  wire                          ena,
  input  wire                          enb,
  input  wire [ADDR_WIDTH_A-1:0]       addra,
  input  wire [ADDR_WIDTH_B-1:0]       addrb,
  input  wire                          wea,
  input  wire [WRITE_DATA_WIDTH_A-1:0] dina,
  output reg  [READ_DATA_WIDTH_B-1:0]  doutb,
  input  wire                          regceb,
  input  wire                          rstb
);
  localparam integer DEPTH = (1 << ADDR_WIDTH_A);

  reg [WRITE_DATA_WIDTH_A-1:0] mem [0:DEPTH-1];

  // Port A: Write
  always @(posedge clka) begin
    if (ena && wea)
      mem[addra] <= dina;
  end

  // Port B: Read (read_first semantics)
  generate
    if (READ_LATENCY_B == 1) begin : g_rl1
      // 1-cycle latency: register mem[addrb] directly to doutb
      always @(posedge clkb) begin
        if (rstb) begin
          doutb <= {READ_DATA_WIDTH_B{1'b0}};
        end else if (enb && regceb) begin
          // For common-clock same-address collision, this samples "old" data
          doutb <= mem[addrb];
        end
      end
    end else begin : g_rlN
      // N-cycle latency (N>=2): pipeline depth = N-1 ahead of doutb
      reg [READ_DATA_WIDTH_B-1:0] pipe [0:READ_LATENCY_B-2];
      integer i;
      always @(posedge clkb) begin
        if (rstb) begin
          for (i = 0; i < READ_LATENCY_B-1; i = i + 1)
            pipe[i] <= {READ_DATA_WIDTH_B{1'b0}};
          doutb <= {READ_DATA_WIDTH_B{1'b0}};
        end else if (enb && regceb) begin
          pipe[0] <= mem[addrb];               // sample current mem value
          for (i = 1; i < READ_LATENCY_B-1; i = i + 1)
            pipe[i] <= pipe[i-1];
          doutb <= pipe[READ_LATENCY_B-2];     // exactly N cycles latency
        end
      end
    end
  endgenerate
endmodule
